magic
tech min2
timestamp 1681500163
<< nwell >>
rect -95 -279 -69 -256
rect -59 -279 -33 -254
rect -23 -279 3 -254
<< ntransistor >>
rect -83 -293 -80 -285
rect -47 -293 -44 -285
rect -11 -293 -8 -285
<< ptransistor >>
rect -83 -273 -80 -265
rect -47 -273 -44 -265
rect -11 -273 -8 -265
<< ndiffusion >>
rect -85 -293 -83 -285
rect -80 -293 -78 -285
rect -49 -293 -47 -285
rect -44 -293 -42 -285
rect -13 -293 -11 -285
rect -8 -293 -6 -285
<< pdiffusion >>
rect -85 -273 -83 -265
rect -80 -273 -78 -265
rect -49 -273 -47 -265
rect -44 -273 -42 -265
rect -13 -273 -11 -265
rect -8 -273 -6 -265
<< ndcontact >>
rect -89 -293 -85 -285
rect -78 -293 -74 -285
rect -53 -293 -49 -285
rect -42 -293 -38 -285
rect -17 -293 -13 -285
rect -6 -293 -2 -285
<< pdcontact >>
rect -89 -273 -85 -265
rect -78 -273 -74 -265
rect -53 -273 -49 -265
rect -42 -273 -38 -265
rect -17 -273 -13 -265
rect -6 -273 -2 -265
<< polysilicon >>
rect -99 -277 -95 -260
rect -83 -265 -80 -262
rect -61 -265 -57 -253
rect -47 -265 -44 -262
rect -11 -265 -8 -260
rect -83 -277 -80 -273
rect -47 -277 -44 -273
rect -11 -276 -8 -273
rect -99 -281 -80 -277
rect -49 -281 -44 -277
rect -83 -285 -80 -281
rect -47 -285 -44 -281
rect -11 -285 -8 -282
rect -83 -296 -80 -293
rect -47 -296 -44 -293
rect -30 -307 -26 -293
rect -11 -298 -8 -293
<< polycontact >>
rect -61 -253 -57 -249
rect -99 -260 -95 -256
rect -11 -260 -8 -256
rect -61 -269 -57 -265
rect -52 -281 -49 -277
rect -30 -293 -26 -289
rect -11 -302 -8 -298
rect -30 -311 -26 -307
<< metal1 >>
rect -99 -256 -95 -252
rect -57 -253 7 -249
rect -95 -260 -11 -256
rect -53 -265 -49 -260
rect -118 -273 -89 -265
rect -118 -330 -113 -273
rect -78 -277 -74 -273
rect -61 -277 -57 -269
rect -42 -277 -38 -273
rect -17 -277 -13 -273
rect -78 -281 -67 -277
rect -61 -281 -52 -277
rect -42 -281 -13 -277
rect -78 -285 -74 -281
rect -106 -293 -89 -285
rect -71 -298 -67 -281
rect -42 -285 -38 -281
rect -30 -289 -26 -281
rect -17 -285 -13 -281
rect -6 -277 -2 -273
rect 3 -277 7 -253
rect -6 -281 7 -277
rect -6 -285 -2 -281
rect -53 -298 -49 -293
rect -71 -302 -11 -298
rect -30 -317 -26 -311
rect 3 -361 7 -281
rect -126 -448 -121 -438
use VCO  VCO_0
timestamp 1680681348
transform 1 0 -148 0 1 -350
box -7 -107 159 29
<< labels >>
rlabel metal1 -28 -315 -28 -315 1 Xor_out
rlabel metal1 5 -279 5 -279 7 VinB
rlabel metal1 -104 -290 -104 -290 3 Gnd
rlabel metal1 -104 -269 -104 -269 3 Vdd
rlabel metal1 -97 -254 -97 -254 5 Vin
rlabel metal1 -123 -446 -123 -446 1 Gnd
<< end >>
