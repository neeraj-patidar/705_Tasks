magic
tech scmos
timestamp 1679443135
<< nwell >>
rect -29 12 66 68
<< polysilicon >>
rect -10 44 -5 47
rect -10 27 -5 39
rect 32 35 37 39
rect -10 6 -5 22
rect 32 16 37 30
rect -10 -10 -5 1
rect 32 -2 37 11
rect 32 -11 37 -7
rect -10 -18 -5 -15
<< ndiffusion >>
rect -15 1 -10 6
rect -5 1 0 6
rect 27 -7 32 -2
rect 37 -7 42 -2
rect -15 -15 -10 -10
rect -5 -15 0 -10
<< pdiffusion >>
rect -15 39 -10 44
rect -5 39 0 44
rect 27 30 32 35
rect 37 30 42 35
rect -15 22 -10 27
rect -5 22 0 27
<< metal1 >>
rect -25 54 -20 64
rect -15 54 0 64
rect 5 54 20 64
rect 25 54 40 64
rect 45 54 59 64
rect -20 44 -15 54
rect 0 35 5 39
rect -20 30 22 35
rect 47 30 52 35
rect -20 27 -15 30
rect 0 16 5 22
rect 0 11 32 16
rect 37 11 43 16
rect 0 6 5 11
rect -20 -2 -15 1
rect -20 -7 22 -2
rect 47 -7 52 -2
rect 0 -10 5 -7
rect -20 -25 -15 -15
rect -25 -35 -20 -25
rect -15 -35 0 -25
rect 5 -35 20 -25
rect 25 -35 40 -25
rect 45 -35 59 -25
<< ntransistor >>
rect -10 1 -5 6
rect 32 -7 37 -2
rect -10 -15 -5 -10
<< ptransistor >>
rect -10 39 -5 44
rect 32 30 37 35
rect -10 22 -5 27
<< polycontact >>
rect 32 11 37 16
<< ndcontact >>
rect -20 1 -15 6
rect 0 1 5 6
rect 22 -7 27 -2
rect 42 -7 47 -2
rect -20 -15 -15 -10
rect 0 -15 5 -10
<< pdcontact >>
rect -20 39 -15 44
rect 0 39 5 44
rect 22 30 27 35
rect 42 30 47 35
rect -20 22 -15 27
rect 0 22 5 27
<< psubstratepcontact >>
rect -20 -35 -15 -25
rect 0 -35 5 -25
rect 20 -35 25 -25
rect 40 -35 45 -25
<< nsubstratencontact >>
rect -20 54 -15 64
rect 0 54 5 64
rect 20 54 25 64
rect 40 54 45 64
<< labels >>
rlabel metal1 12 60 12 60 1 Vdd
rlabel metal1 50 -5 50 -5 1 Vdd
rlabel metal1 13 -31 13 -31 1 Gnd
rlabel metal1 50 32 50 32 1 Gnd
rlabel polysilicon -7 10 -7 10 1 Vin
rlabel metal1 40 14 40 14 1 Vout
<< end >>
